`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/17/2020 09:48:57 PM
// Design Name: 
// Module Name: Controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Controller(instruction, funct, 
                  regDst, ALUSource, MemToReg, regWrite, MemRead, MemWrite, Jump, BranchJump, ALUOp, MulOp, MemDataType);
    input [5:0] instruction, funct;
    output reg [1:0] MemDataType;
    output reg regDst, ALUSource, MemToReg, regWrite, MemRead, MemWrite, MulOp, Jump;
    output reg [2:0] BranchJump;
    output reg [4:0] ALUOp;
    
    initial begin
        MulOp <= 0;
        MemDataType <= 0;
        regDst <= 0;
        ALUSource <= 0;
        MemToReg <= 0;
        regWrite <= 0;
        MemRead <= 0;
        MemWrite <= 0;
        Jump <= 0;
        BranchJump <= 3'b0;
        ALUOp <= 5'b0;
    end
    
    always @ (*) begin
        MulOp <= 0;
        MemDataType <= 0;
        regDst <= 0;
        ALUSource <= 0;
        MemToReg <= 0;
        regWrite <= 0;
        MemRead <= 0;
        MemWrite <= 0;
        Jump <= 0;
        BranchJump <= 3'b0;
        ALUOp <= 5'b0;
    
        case (instruction)
            6'b000000: begin // r-type
                regDst <= 1'b0;
                ALUSource <= 1'b0;
                MemToReg <= 1'b1;
                regWrite <= 1'b1;
                MemRead <= 1'b0;
                MemWrite <= 1'b0;
                BranchJump <= 3'b000;
                ALUOp <= 5'b00000;
                case (funct) 
                    6'b011000: MulOp <= 1;
                    6'b011001: MulOp <= 1;
                    default: MulOp <= 0;
                endcase
            end
            6'b001000: begin // addi
                  regDst <= 1;
                  ALUSource <= 1;
                  MemToReg <= 1;
                  regWrite <= 1;
                  MemRead <= 0;
                  MemWrite <= 0;
                  BranchJump <= 0;
                  ALUOp <= 5'b00010; //  add Code
                  MulOp <= 0;
            end
            6'b001001: begin // addiu
                regDst <= 1;
                ALUSource <= 1;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00111; // todo: Change to addu Code
                MulOp <= 0;
            end
            6'b011100: begin // special2  madd/msub
                regDst <= 0;
                ALUSource <= 0;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b01000; // 
                MulOp <= 1;
            end
            6'b011111: begin // special3  seb/seh
                regDst <= 0;
                ALUSource <= 0;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b01001; // 
                MulOp <= 0;
            end
            6'b100011: begin // lw
                MemDataType <= 2'b10;
                regDst <= 1;
                ALUSource <= 1;
                MemToReg <= 0;
                regWrite <= 1;
                MemRead <= 1;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00010; // add Code
                MulOp <= 0;
            end
            6'b101011: begin // sw
                MemDataType <= 2'b10;
                ALUSource <= 1;
                regWrite <= 0;
                MemRead <= 0;
                MemWrite <= 1;
                BranchJump <= 0;
                ALUOp <= 5'b00010; // add Code
                MulOp <= 0;
            end
            6'b100000: begin // lb
                MemDataType <= 2'b00;
                regDst <= 0;
                ALUSource <= 1;
                MemToReg <= 0;
                regWrite <= 1;
                MemRead <= 1;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00010; // add Code
                MulOp <= 0;
            end
            6'b100001: begin //lh
                MemDataType <= 2'b01;
                regDst <= 0;
                ALUSource <= 1;
                MemToReg <= 0;
                regWrite <= 1;
                MemRead <= 1;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00010; // add Code
                MulOp <= 0;
            end
            6'b101000: begin // sb
                MemDataType <= 2'b00;
                ALUSource <= 1;
                regWrite <= 0;
                MemRead <= 0;
                MemWrite <= 1;
                BranchJump <= 0;
                ALUOp <= 5'b00010; // add Code
                MulOp <= 0;
            end
            6'b101001: begin // sh
                MemDataType <= 2'b01;
                ALUSource <= 1;
                regWrite <= 0;
                MemRead <= 0;
                MemWrite <= 1;
                BranchJump <= 0;
                ALUOp <= 5'b00010; // add Code
                MulOp <= 0;
            end
            6'b001111: begin // lui
                MemDataType <= 2'b00;
                regDst <= 1;   // 1 for rt, 0 for rd
                ALUSource <= 1; // 1 for offset, 0 for readdata2
                MemToReg <= 1; // 1 for alu output, 0 for datamemory output
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b10100; // lui Code
                MulOp <= 0;
            end
            6'b000001: begin // bltz/ bgez
                Jump <= 1;
                BranchJump <= 3'b100;
                ALUOp <= 5'b00110; // todo: Change to sub Code
            end
            6'b000100: begin // beq
                Jump <= 1;
                BranchJump <= 3'b001;
                ALUOp <= 5'b00110; // sub Code
            end
            6'b000101: begin // bne
                Jump <= 1;
                BranchJump <= 3'b010;
                ALUOp <= 5'b00110; // sub Code
                MulOp <= 0;
            end
            6'b000111: begin // bgtz
                Jump <= 1;
                BranchJump <= 3'b101;
                ALUOp <= 5'b00110; // todo: Change to sub Code
            end
            6'b000110: begin // blez
                Jump <= 1;
                BranchJump <= 3'b110;
                ALUOp <= 5'b00110; // todo: Change to sub Code
            end
            6'b000010: begin // j // reqires datapath modification
                Jump <= 1;
                BranchJump <= 3'b011;
                ALUOp <= 5'b00110; // todo: Change to sub Code
            end
            6'b000011: begin // jal
                Jump <= 1;
                BranchJump <= 3'b011;
                ALUOp <= 5'b00110; // todo: Change to sub Code
            end
            6'b001100: begin // andi
                regDst <= 1;
                ALUSource <= 1;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00001; // change to and code
                MulOp <= 0;
            end
            6'b001101: begin // ori
                regDst <= 1;
                ALUSource <= 1;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00011; // change to or code
                MulOp <= 0;
            end
            6'b001110: begin // xori
                regDst <= 1;
                ALUSource <= 1;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00100; // change to xor code
                MulOp <= 0;
            end
            6'b001010: begin // slti
                regDst <= 1;
                ALUSource <= 1;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b00101; // change to slt code
                MulOp <= 0;
            end
            6'b001011: begin // sltiu
                regDst <= 1;
                ALUSource <= 1;
                MemToReg <= 1;
                regWrite <= 1;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 0;
                ALUOp <= 5'b01011; // change to sltu code
                MulOp <= 0;
            end
            default: begin
                MulOp <= 0;
                MemDataType <= 0;
                regDst <= 0;
                ALUSource <= 0;
                MemToReg <= 0;
                regWrite <= 0;
                MemRead <= 0;
                MemWrite <= 0;
                BranchJump <= 3'b0;
                ALUOp <= 5'b0;
            end 
        endcase
    end
endmodule